`timescale 1ns / 1ps

module andGate
    (
    input  a,b,
    output c
    );
    
    assign c = a & b;
    
endmodule
